LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY part5 IS
		PORT ( SW : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
		HEX0 : OUT STD_LOGIC_VECTOR(0 TO 6);
		HEX1 : OUT STD_LOGIC_VECTOR(0 TO 6);
		HEX2 : OUT STD_LOGIC_VECTOR(0 TO 6);
		HEX3 : OUT STD_LOGIC_VECTOR(0 TO 6);
		HEX4 : OUT STD_LOGIC_VECTOR(0 TO 6));
END part5;

ARCHITECTURE Behavior OF part5 IS
	
	COMPONENT mux_3bit_5to1
		PORT ( S, U, V, W, X, Y : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		M : OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
	END COMPONENT;

	COMPONENT char_7seg
		PORT ( C : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		Display : OUT STD_LOGIC_VECTOR(0 TO 6));
	END COMPONENT;

	SIGNAL M, N, O, P, Q : STD_LOGIC_VECTOR(2 DOWNTO 0);
	
	BEGIN
	M0: mux_3bit_5to1 PORT MAP (SW(17 DOWNTO 15), SW(14 DOWNTO 12), SW(11 DOWNTO 9), SW(8 DOWNTO 6), SW(5 DOWNTO 3), SW(2 DOWNTO 0), M);
	H0: char_7seg PORT MAP (M, HEX0);

	M1: mux_3bit_5to1 PORT MAP (SW(17 DOWNTO 15), SW(11 DOWNTO 9), SW(8 DOWNTO 6), SW(5 DOWNTO 3), SW(2 DOWNTO 0), SW(14 DOWNTO 12), N);
	H1: char_7seg PORT MAP (N, HEX1);

	M2: mux_3bit_5to1 PORT MAP (SW(17 DOWNTO 15), SW(8 DOWNTO 6), SW(5 DOWNTO 3), SW(2 DOWNTO 0), SW(14 DOWNTO 12), SW(11 DOWNTO 9), O);
	H2: char_7seg PORT MAP (O, HEX2);

	M3: mux_3bit_5to1 PORT MAP (SW(17 DOWNTO 15), SW(5 DOWNTO 3), SW(2 DOWNTO 0), SW(14 DOWNTO 12), SW(11 DOWNTO 9), SW(8 DOWNTO 6), P);
	H3: char_7seg PORT MAP (P, HEX3);

	M4: mux_3bit_5to1 PORT MAP (SW(17 DOWNTO 15), SW(2 DOWNTO 0), SW(14 DOWNTO 12), SW(11 DOWNTO 9), SW(8 DOWNTO 6), SW(5 DOWNTO 3), Q);
	H4: char_7seg PORT MAP (Q, HEX4);

END Behavior;