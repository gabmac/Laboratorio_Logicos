LIBRARY ieee;
USE ieee.std_logic_1164.all;
ENTITY P5 IS
PORT ( 
	SW : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	KEY :IN STD_LOGIC_VECTOR(1 DOWNTO 0);
	HEX0,HEX1,HEX2,HEX3,HEX4,HEX5,HEX6,HEX7:OUT STD_LOGIC_VECTOR(0 TO 6));
END P5;
	ARCHITECTURE Structural OF P5 IS
	COMPONENT FLIPFLOP IS
	PORT ( 
	CLK,D, RESET : IN STD_LOGIC;
	Q : OUT STD_LOGIC);
END COMPONENT;

	COMPONENT Parte5 IS
	PORT (  SW : IN std_logic_vector (3 DOWNTO 0) ;
	HEX0 : OUT std_logic_vector (0 TO 6)  ) ;
END COMPONENT;
	
	SIGNAL VECTOR: STD_LOGIC_VECTOR(15 DOWNTO 0);
	
BEGIN
	-- Valor Atual --
	P0: Parte5 PORT MAP(SW(3 DOWNTO 0),HEX4);
	P1: Parte5 PORT MAP(SW(7 DOWNTO 4),HEX5);
	P2: Parte5 PORT MAP(SW(11 DOWNTO 8),HEX6);
	P3: Parte5 PORT MAP(SW(15 DOWNTO 12),HEX7);
	
	-- Memoriza --
	
	FF0: FLIPFLOP PORT MAP (KEY(0),SW(0),KEY(1),VECTOR(0));
	FF1: FLIPFLOP PORT MAP (KEY(0),SW(1),KEY(1),VECTOR(1));
	FF2: FLIPFLOP PORT MAP (KEY(0),SW(2),KEY(1),VECTOR(2));
	FF3: FLIPFLOP PORT MAP (KEY(0),SW(3),KEY(1),VECTOR(3));
	FF4: FLIPFLOP PORT MAP (KEY(0),SW(4),KEY(1),VECTOR(4));
	FF5: FLIPFLOP PORT MAP (KEY(0),SW(5),KEY(1),VECTOR(5));
	FF6: FLIPFLOP PORT MAP (KEY(0),SW(6),KEY(1),VECTOR(6));
	FF7: FLIPFLOP PORT MAP (KEY(0),SW(7),KEY(1),VECTOR(7));
	FF8: FLIPFLOP PORT MAP (KEY(0),SW(8),KEY(1),VECTOR(8));
	FF9: FLIPFLOP PORT MAP (KEY(0),SW(9),KEY(1),VECTOR(9));
	FF10: FLIPFLOP PORT MAP (KEY(0),SW(10),KEY(1),VECTOR(10));
	FF11: FLIPFLOP PORT MAP (KEY(0),SW(11),KEY(1),VECTOR(11));
	FF12: FLIPFLOP PORT MAP (KEY(0),SW(12),KEY(1),VECTOR(12));
	FF13: FLIPFLOP PORT MAP (KEY(0),SW(13),KEY(1),VECTOR(13));
	FF14: FLIPFLOP PORT MAP (KEY(0),SW(14),KEY(1),VECTOR(14));
	FF15: FLIPFLOP PORT MAP (KEY(0),SW(15),KEY(1),VECTOR(15));
	
	P4: Parte5 PORT MAP(VECTOR(3 DOWNTO 0),HEX0);
	P5: Parte5 PORT MAP(VECTOR(7 DOWNTO 4),HEX1);
	P6: Parte5 PORT MAP(VECTOR(11 DOWNTO 8),HEX2);
	P7: Parte5 PORT MAP(VECTOR(15 DOWNTO 12),HEX3);
	
END Structural;