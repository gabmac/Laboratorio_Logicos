LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Exp1b IS
	PORT ( SW : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
	LEDR : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
	LEDG : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END Exp1b;

ARCHITECTURE Behavior OF Exp1b IS
	BEGIN
	LEDR <= SW;
	LEDG(0) <= (NOT (SW(17)) AND SW(0)) OR (SW(17) AND SW(8));
	LEDG(1) <= (NOT (SW(17)) AND SW(1)) OR (SW(17) AND SW(9));
	LEDG(2) <= (NOT (SW(17)) AND SW(2)) OR (SW(17) AND SW(10));
	LEDG(3) <= (NOT (SW(17)) AND SW(3)) OR (SW(17) AND SW(11));
	LEDG(4) <= (NOT (SW(17)) AND SW(4)) OR (SW(17) AND SW(12));
	LEDG(5) <= (NOT (SW(17)) AND SW(5)) OR (SW(17) AND SW(13));
	LEDG(6) <= (NOT (SW(17)) AND SW(6)) OR (SW(17) AND SW(14));
	LEDG(7) <= (NOT (SW(17)) AND SW(7)) OR (SW(17) AND SW(15));
END Behavior;
