LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Lab2D IS
	PORT ( SW : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
	HEX0, HEX1, HEX6, HEX4 : OUT STD_LOGIC_VECTOR(0 TO 6);
	LEDR, LEDG : OUT STD_LOGIC_VECTOR(8 DOWNTO 0));
	 
END Lab2D;

ARCHITECTURE Behavior OF Lab2D IS
		
		COMPONENT DISP
		PORT ( SW : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	Display : OUT STD_LOGIC_VECTOR(0 TO 6));
	END COMPONENT;
	
	COMPONENT Somador IS
	PORT (Cin : IN STD_LOGIC;
	Saida : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
	Entrada : IN STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

	COMPONENT Tradutor IS
		PORT (V : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		C, O: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
	END COMPONENT;
		
		SIGNAL S: STD_LOGIC_VECTOR(4 DOWNTO 0);
		SIGNAL D, U : STD_LOGIC_VECTOR(3 DOWNTO 0);
		
		BEGIN
		
	LEDR <= SW;
	
	H6: DISP PORT MAP(SW(7 DOWNTO 4),HEX6);
	H4: DISP PORT MAP(SW(3 DOWNTO 0),HEX4);
	
	LEDG(8) <= ((SW(7) AND (SW(6) OR SW(5))) OR (SW(3) AND (SW(2) OR SW(1))));
	
	SOMA:  Somador PORT MAP(SW(8),S,SW(7 DOWNTO 0));
	
	T: Tradutor PORT MAP(S, D, U);
	
	
	H1: DISP PORT MAP(D,HEX1);
	H0: DISP PORT MAP(U,HEX0);
	
	
	
END BEHAVIOR;