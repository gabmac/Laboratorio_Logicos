LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Exp2a IS
	PORT ( SW : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
	LEDR : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
	HEX0 : OUT STD_LOGIC_VECTOR(0 TO 6);
	HEX1 : OUT STD_LOGIC_VECTOR(0 TO 6);
	HEX2 : OUT STD_LOGIC_VECTOR(0 TO 6);
	HEX3 : OUT STD_LOGIC_VECTOR(0 TO 6));
END Exp2a;

ARCHITECTURE Behavior OF Exp2a IS
	
	COMPONENT Exp1d
		PORT ( SW : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		Display : OUT STD_LOGIC_VECTOR(0 TO 6));
	END COMPONENT;


	BEGIN
	LEDR <= SW;
	
	H0: Exp1d PORT MAP (SW(3 DOWNTO 0), HEX0);
	H1: Exp1d PORT MAP (SW(7 DOWNTO 4), HEX1);
	H2: Exp1d PORT MAP (SW(11 DOWNTO 8), HEX2);
	H3: Exp1d PORT MAP (SW(15 DOWNTO 12), HEX3);
	
END Behavior;
 	