--		Julio Alves Mesquita da Silva			156061 	--
--		Gabriel Bonani Machado					155416	--

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
ENTITY Main IS
PORT ( 
	CLOCK_50: IN STD_LOGIC;
	SW: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
	HEX0:OUT STD_LOGIC_VECTOR(0 TO 6));
END Main;
	ARCHITECTURE Structural OF Main IS
	
	
	Component seg IS
	PORT (  SW : IN std_logic_vector (3 DOWNTO 0) ;
	HEX0 : OUT std_logic_vector (0 TO 6)  ) ;
END COMPONENT;

	
	SIGNAL C: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
	SIGNAL Estado : std_logic_vector(28 DOWNTO 0) := "00000000000000000000000000000";
	
BEGIN
	
	PROCESS(Estado)

  BEGIN	
	 
    IF ( rising_edge(CLOCK_50)) THEN
      Estado <= Estado + '1';

    END IF;
	 

	IF(Estado =  "11101110011010110010100000000") THEN
		Estado <= "00000000000000000000000000000";
	END IF;
		
	IF ((Estado > "00000000000000000000000000000") AND (Estado < "00010111110101111000010000000")) THEN
		C <= 	 "0000";
	ELSIF ((Estado > "00010111110101111000010000000") AND (Estado < "00101111101011110000100000000")) THEN
		C <= 	 "0001";
	ELSIF ((Estado > "00101111101011110000100000000") AND (Estado < "01000111100001101000110000000")) THEN
		C <= 	 "0010";
	ELSIF ((Estado > "01000111100001101000110000000") AND (Estado < "01011111010111100001000000000")) THEN
		C <= 	 "0011";
	ELSIF ((Estado > "01011111010111100001000000000") AND (Estado < "01110111001101011001010000000")) THEN
		C <= 	 "0100";
	ELSIF ((Estado > "01110111001101011001010000000") AND (Estado < "10001111000011010001100000000")) THEN
		C <= 	 "0101";
	ELSIF ((Estado > "10001111000011010001100000000") AND (Estado < "10100110111001001001110000000")) THEN
		C <= 	 "0110";
	ELSIF ((Estado > "10100110111001001001110000000") AND (Estado < "10111110101111000010000000000")) THEN
		C <= 	 "0111";
	ELSIF ((Estado > "10111110101111000010000000000") AND (Estado < "11010110100100111010010000000")) THEN
		C <= 	 "1000";
	ELSIF ((Estado > "11010110100100111010010000000")) THEN
		C <= 	 "1001";
	ELSE C <= C;
	END IF;
			
	END PROCESS;
	
			
	
	H0: seg PORT MAP(C, HEX0);

	
END Structural;